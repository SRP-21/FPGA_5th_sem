`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 26.12.2025 22:23:02
// Design Name: 
// Module Name: state_predictor
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module state_predictor (

    input  signed [15:0] X0, X1,X2,X3,X4,X5,

    input  signed [15:0]
        P0,  P1,  P2,  P3,  P4,  P5,
        P6,  P7,  P8,  P9,  P10, P11,
        P12, P13, P14, P15, P16, P17,
        P18, P19, P20, P21, P22, P23,
        P24, P25, P26, P27, P28, P29,
        P30, P31, P32, P33, P34, P35,

    output reg signed [31:0] Xn0, Xn1,Xn2,Xn3,Xn4,Xn5,

   output reg signed [31:0]
        Pn0,  Pn1,  Pn2,  Pn3,  Pn4,  Pn5,
        Pn6,  Pn7,  Pn8,  Pn9,  Pn10, Pn11,
        Pn12, Pn13, Pn14, Pn15, Pn16, Pn17,
        Pn18, Pn19, Pn20, Pn21, Pn22, Pn23,
        Pn24, Pn25, Pn26, Pn27, Pn28, Pn29,
        Pn30, Pn31, Pn32, Pn33, Pn34, Pn35
);


wire signed [15:0] F [0:35];
wire signed [15:0] Q [0:35];



 parameter signed [15:0] ONE  = 16'sd1;
 parameter signed [15:0] ZERO = 16'sd0;
 parameter signed [15:0] Dt   = 16'sd1;
 parameter signed [15:0] CovP = 16'sd1;
 parameter signed [15:0] CovV = 16'sd10;

assign F0  = ONE;   assign F1  = ZERO; assign F2  = ZERO; assign F3  = Dt;    assign F4  = ZERO; assign F5  = ZERO;
assign F6  = ZERO;  assign F7  = ONE;  assign F8  = ZERO; assign F9  = ZERO;  assign F10 = Dt;   assign F11 = ZERO;
assign F12 = ZERO;  assign F13 = ZERO; assign F14 = ONE; assign F15 = ZERO;  assign F16 = ZERO; assign F17 = Dt;
assign F18 = ZERO;  assign F19 = ZERO; assign F20 = ZERO; assign F21 = ONE;   assign F22 = ZERO; assign F23 = ZERO;
assign F24 = ZERO;  assign F25 = ZERO; assign F26 = ZERO; assign F27 = ZERO;  assign F28 = ONE;  assign F29 = ZERO;
assign F30 = ZERO;  assign F31 = ZERO; assign F32 = ZERO; assign F33 = ZERO;  assign F34 = ZERO; assign F35 = ONE;

assign Q0 = CovP; assign Q1 = ZERO; assign Q2 = ZERO; assign Q3 = ZERO; assign Q4 = ZERO; assign Q5 = ZERO;
assign Q6 = ZERO; assign Q7 = CovV; assign Q8 = ZERO; assign Q9 = ZERO; assign Q10 = ZERO; assign Q11 = ZERO;
assign Q12 = ZERO; assign Q13 = ZERO; assign Q14 = CovP; assign Q15 = ZERO; assign Q16 = ZERO; assign Q17 = ZERO;
assign Q18 = ZERO; assign Q19 = ZERO; assign Q20 = ZERO; assign Q21 = CovV; assign Q22 = ZERO; assign Q23 = ZERO;
assign Q24 = ZERO; assign Q25 = ZERO; assign Q26 = ZERO; assign Q27 = ZERO; assign Q28 = CovP; assign Q29 = ZERO;
assign Q30 = ZERO; assign Q31 = ZERO; assign Q32 = ZERO; assign Q33 = ZERO; assign Q34 = CovP; assign Q35 = CovV;

always @(*) begin
 Xn0 = F0*X0 + F1*X1 + F2*X2 + F3*X3 + F4*X4 + F5*X5;
 Xn1 = F6*X0 + F7*X1 + F8*X2 + F9*X3 + F10*X4 + F11*X5;
 Xn2 = F12*X0 + F13*X1 + F14*X2 + F15*X3 + F16*X4 + F17*X5;
 Xn3 = F18*X0 + F19*X1 + F20*X2 + F21*X3 + F22*X4 + F23*X5;
 Xn4 = F24*X0 + F25*X1 + F26*X2 + F27*X3 + F28*X4 + F29*X5;
 Xn5 = F30*X0 + F31*X1 + F32*X2 + F33*X3 + F34*X4 + F35*X5;

 Pn0 = (F0*P0 + F0*P1 + F0*P2 + F0*P3 + F0*P4 + F0*P5)*F5 + 
    (F1*P6 + F1*P7 + F1*P8 + F1*P9 + F1*P10 + F1*P11)*F5 + 
    (F2*P12 + F2*P13 + F2*P14 + F2*P15 + F2*P16 + F2*P17)*F5 + 
    (F3*P18 + F3*P19 + F3*P20 + F3*P21 + F3*P22 + F3*P23)*F5 + 
    (F4*P24 + F4*P25 + F4*P26 + F4*P27 + F4*P28 + F4*P29)*F5 + 
    (F5*P30 + F5*P31 + F5*P32 + F5*P33 + F5*P34 + F5*P35)*F5 + Q0;

 Pn1 = (F0*P0 + F0*P1 + F0*P2 + F0*P3 + F0*P4 + F0*P5)*F11 + 
    (F1*P6 + F1*P7 + F1*P8 + F1*P9 + F1*P10 + F1*P11)*F11 + 
    (F2*P12 + F2*P13 + F2*P14 + F2*P15 + F2*P16 + F2*P17)*F11 + 
    (F3*P18 + F3*P19 + F3*P20 + F3*P21 + F3*P22 + F3*P23)*F11 + 
    (F4*P24 + F4*P25 + F4*P26 + F4*P27 + F4*P28 + F4*P29)*F11 + 
    (F5*P30 + F5*P31 + F5*P32 + F5*P33 + F5*P34 + F5*P35)*F11 + Q1;

 Pn2 = (F0*P0 + F0*P1 + F0*P2 + F0*P3 + F0*P4 + F0*P5)*F17 + 
    (F1*P6 + F1*P7 + F1*P8 + F1*P9 + F1*P10 + F1*P11)*F17 + 
    (F2*P12 + F2*P13 + F2*P14 + F2*P15 + F2*P16 + F2*P17)*F17 + 
    (F3*P18 + F3*P19 + F3*P20 + F3*P21 + F3*P22 + F3*P23)*F17 + 
    (F4*P24 + F4*P25 + F4*P26 + F4*P27 + F4*P28 + F4*P29)*F17 + 
    (F5*P30 + F5*P31 + F5*P32 + F5*P33 + F5*P34 + F5*P35)*F17 + Q2;

 Pn3 = (F0*P0 + F0*P1 + F0*P2 + F0*P3 + F0*P4 + F0*P5)*F23 + 
    (F1*P6 + F1*P7 + F1*P8 + F1*P9 + F1*P10 + F1*P11)*F23 + 
    (F2*P12 + F2*P13 + F2*P14 + F2*P15 + F2*P16 + F2*P17)*F23 + 
    (F3*P18 + F3*P19 + F3*P20 + F3*P21 + F3*P22 + F3*P23)*F23 + 
    (F4*P24 + F4*P25 + F4*P26 + F4*P27 + F4*P28 + F4*P29)*F23 + 
    (F5*P30 + F5*P31 + F5*P32 + F5*P33 + F5*P34 + F5*P35)*F23 + Q3;

 Pn4 = (F0*P0 + F0*P1 + F0*P2 + F0*P3 + F0*P4 + F0*P5)*F29 + 
    (F1*P6 + F1*P7 + F1*P8 + F1*P9 + F1*P10 + F1*P11)*F29 + 
    (F2*P12 + F2*P13 + F2*P14 + F2*P15 + F2*P16 + F2*P17)*F29 + 
    (F3*P18 + F3*P19 + F3*P20 + F3*P21 + F3*P22 + F3*P23)*F29 + 
    (F4*P24 + F4*P25 + F4*P26 + F4*P27 + F4*P28 + F4*P29)*F29 + 
    (F5*P30 + F5*P31 + F5*P32 + F5*P33 + F5*P34 + F5*P35)*F29 + Q4;

 Pn5 = (F0*P0 + F0*P1 + F0*P2 + F0*P3 + F0*P4 + F0*P5)*F35 + 
    (F1*P6 + F1*P7 + F1*P8 + F1*P9 + F1*P10 + F1*P11)*F35 + 
    (F2*P12 + F2*P13 + F2*P14 + F2*P15 + F2*P16 + F2*P17)*F35 + 
    (F3*P18 + F3*P19 + F3*P20 + F3*P21 + F3*P22 + F3*P23)*F35 + 
    (F4*P24 + F4*P25 + F4*P26 + F4*P27 + F4*P28 + F4*P29)*F35 + 
    (F5*P30 + F5*P31 + F5*P32 + F5*P33 + F5*P34 + F5*P35)*F35 + Q5;

 Pn6 = (F6*P0 + F6*P1 + F6*P2 + F6*P3 + F6*P4 + F6*P5)*F5 + 
    (F7*P6 + F7*P7 + F7*P8 + F7*P9 + F7*P10 + F7*P11)*F5 + 
    (F8*P12 + F8*P13 + F8*P14 + F8*P15 + F8*P16 + F8*P17)*F5 + 
    (F9*P18 + F9*P19 + F9*P20 + F9*P21 + F9*P22 + F9*P23)*F5 + 
    (F10*P24 + F10*P25 + F10*P26 + F10*P27 + F10*P28 + F10*P29)*F5 + 
    (F11*P30 + F11*P31 + F11*P32 + F11*P33 + F11*P34 + F11*P35)*F5 + Q6;

 Pn7 = (F6*P0 + F6*P1 + F6*P2 + F6*P3 + F6*P4 + F6*P5)*F11 + 
    (F7*P6 + F7*P7 + F7*P8 + F7*P9 + F7*P10 + F7*P11)*F11 + 
    (F8*P12 + F8*P13 + F8*P14 + F8*P15 + F8*P16 + F8*P17)*F11 + 
    (F9*P18 + F9*P19 + F9*P20 + F9*P21 + F9*P22 + F9*P23)*F11 + 
    (F10*P24 + F10*P25 + F10*P26 + F10*P27 + F10*P28 + F10*P29)*F11 + 
    (F11*P30 + F11*P31 + F11*P32 + F11*P33 + F11*P34 + F11*P35)*F11 + Q7;

 Pn8 = (F6*P0 + F6*P1 + F6*P2 + F6*P3 + F6*P4 + F6*P5)*F17 + 
    (F7*P6 + F7*P7 + F7*P8 + F7*P9 + F7*P10 + F7*P11)*F17 + 
    (F8*P12 + F8*P13 + F8*P14 + F8*P15 + F8*P16 + F8*P17)*F17 + 
    (F9*P18 + F9*P19 + F9*P20 + F9*P21 + F9*P22 + F9*P23)*F17 + 
    (F10*P24 + F10*P25 + F10*P26 + F10*P27 + F10*P28 + F10*P29)*F17 + 
    (F11*P30 + F11*P31 + F11*P32 + F11*P33 + F11*P34 + F11*P35)*F17 + Q8;

 Pn9 = (F6*P0 + F6*P1 + F6*P2 + F6*P3 + F6*P4 + F6*P5)*F23 + 
    (F7*P6 + F7*P7 + F7*P8 + F7*P9 + F7*P10 + F7*P11)*F23 + 
    (F8*P12 + F8*P13 + F8*P14 + F8*P15 + F8*P16 + F8*P17)*F23 + 
    (F9*P18 + F9*P19 + F9*P20 + F9*P21 + F9*P22 + F9*P23)*F23 + 
    (F10*P24 + F10*P25 + F10*P26 + F10*P27 + F10*P28 + F10*P29)*F23 + 
    (F11*P30 + F11*P31 + F11*P32 + F11*P33 + F11*P34 + F11*P35)*F23 + Q9;

 Pn10 = (F6*P0 + F6*P1 + F6*P2 + F6*P3 + F6*P4 + F6*P5)*F29 + 
    (F7*P6 + F7*P7 + F7*P8 + F7*P9 + F7*P10 + F7*P11)*F29 + 
    (F8*P12 + F8*P13 + F8*P14 + F8*P15 + F8*P16 + F8*P17)*F29 + 
    (F9*P18 + F9*P19 + F9*P20 + F9*P21 + F9*P22 + F9*P23)*F29 + 
    (F10*P24 + F10*P25 + F10*P26 + F10*P27 + F10*P28 + F10*P29)*F29 + 
    (F11*P30 + F11*P31 + F11*P32 + F11*P33 + F11*P34 + F11*P35)*F29 + Q10;

 Pn11 = (F6*P0 + F6*P1 + F6*P2 + F6*P3 + F6*P4 + F6*P5)*F35 + 
    (F7*P6 + F7*P7 + F7*P8 + F7*P9 + F7*P10 + F7*P11)*F35 + 
    (F8*P12 + F8*P13 + F8*P14 + F8*P15 + F8*P16 + F8*P17)*F35 + 
    (F9*P18 + F9*P19 + F9*P20 + F9*P21 + F9*P22 + F9*P23)*F35 + 
    (F10*P24 + F10*P25 + F10*P26 + F10*P27 + F10*P28 + F10*P29)*F35 + 
    (F11*P30 + F11*P31 + F11*P32 + F11*P33 + F11*P34 + F11*P35)*F35 + Q11;

 Pn12 = (F12*P0 + F12*P1 + F12*P2 + F12*P3 + F12*P4 + F12*P5)*F5 + 
    (F13*P6 + F13*P7 + F13*P8 + F13*P9 + F13*P10 + F13*P11)*F5 + 
    (F14*P12 + F14*P13 + F14*P14 + F14*P15 + F14*P16 + F14*P17)*F5 + 
    (F15*P18 + F15*P19 + F15*P20 + F15*P21 + F15*P22 + F15*P23)*F5 + 
    (F16*P24 + F16*P25 + F16*P26 + F16*P27 + F16*P28 + F16*P29)*F5 + 
    (F17*P30 + F17*P31 + F17*P32 + F17*P33 + F17*P34 + F17*P35)*F5 + Q12;

 Pn13 = (F12*P0 + F12*P1 + F12*P2 + F12*P3 + F12*P4 + F12*P5)*F11 + 
    (F13*P6 + F13*P7 + F13*P8 + F13*P9 + F13*P10 + F13*P11)*F11 + 
    (F14*P12 + F14*P13 + F14*P14 + F14*P15 + F14*P16 + F14*P17)*F11 + 
    (F15*P18 + F15*P19 + F15*P20 + F15*P21 + F15*P22 + F15*P23)*F11 + 
    (F16*P24 + F16*P25 + F16*P26 + F16*P27 + F16*P28 + F16*P29)*F11 + 
    (F17*P30 + F17*P31 + F17*P32 + F17*P33 + F17*P34 + F17*P35)*F11 + Q13;

 Pn14 = (F12*P0 + F12*P1 + F12*P2 + F12*P3 + F12*P4 + F12*P5)*F17 + 
    (F13*P6 + F13*P7 + F13*P8 + F13*P9 + F13*P10 + F13*P11)*F17 + 
    (F14*P12 + F14*P13 + F14*P14 + F14*P15 + F14*P16 + F14*P17)*F17 + 
    (F15*P18 + F15*P19 + F15*P20 + F15*P21 + F15*P22 + F15*P23)*F17 + 
    (F16*P24 + F16*P25 + F16*P26 + F16*P27 + F16*P28 + F16*P29)*F17 + 
    (F17*P30 + F17*P31 + F17*P32 + F17*P33 + F17*P34 + F17*P35)*F17 + Q14;

 Pn15 = (F12*P0 + F12*P1 + F12*P2 + F12*P3 + F12*P4 + F12*P5)*F23 + 
    (F13*P6 + F13*P7 + F13*P8 + F13*P9 + F13*P10 + F13*P11)*F23 + 
    (F14*P12 + F14*P13 + F14*P14 + F14*P15 + F14*P16 + F14*P17)*F23 + 
    (F15*P18 + F15*P19 + F15*P20 + F15*P21 + F15*P22 + F15*P23)*F23 + 
    (F16*P24 + F16*P25 + F16*P26 + F16*P27 + F16*P28 + F16*P29)*F23 + 
    (F17*P30 + F17*P31 + F17*P32 + F17*P33 + F17*P34 + F17*P35)*F23 + Q15;

 Pn16 = (F12*P0 + F12*P1 + F12*P2 + F12*P3 + F12*P4 + F12*P5)*F29 + 
    (F13*P6 + F13*P7 + F13*P8 + F13*P9 + F13*P10 + F13*P11)*F29 + 
    (F14*P12 + F14*P13 + F14*P14 + F14*P15 + F14*P16 + F14*P17)*F29 + 
    (F15*P18 + F15*P19 + F15*P20 + F15*P21 + F15*P22 + F15*P23)*F29 + 
    (F16*P24 + F16*P25 + F16*P26 + F16*P27 + F16*P28 + F16*P29)*F29 + 
    (F17*P30 + F17*P31 + F17*P32 + F17*P33 + F17*P34 + F17*P35)*F29 + Q16;

 Pn17 = (F12*P0 + F12*P1 + F12*P2 + F12*P3 + F12*P4 + F12*P5)*F35 + 
    (F13*P6 + F13*P7 + F13*P8 + F13*P9 + F13*P10 + F13*P11)*F35 + 
    (F14*P12 + F14*P13 + F14*P14 + F14*P15 + F14*P16 + F14*P17)*F35 + 
    (F15*P18 + F15*P19 + F15*P20 + F15*P21 + F15*P22 + F15*P23)*F35 + 
    (F16*P24 + F16*P25 + F16*P26 + F16*P27 + F16*P28 + F16*P29)*F35 + 
    (F17*P30 + F17*P31 + F17*P32 + F17*P33 + F17*P34 + F17*P35)*F35 + Q17;

 Pn18 = (F18*P0 + F18*P1 + F18*P2 + F18*P3 + F18*P4 + F18*P5)*F5 + 
    (F19*P6 + F19*P7 + F19*P8 + F19*P9 + F19*P10 + F19*P11)*F5 + 
    (F20*P12 + F20*P13 + F20*P14 + F20*P15 + F20*P16 + F20*P17)*F5 + 
    (F21*P18 + F21*P19 + F21*P20 + F21*P21 + F21*P22 + F21*P23)*F5 + 
    (F22*P24 + F22*P25 + F22*P26 + F22*P27 + F22*P28 + F22*P29)*F5 + 
    (F23*P30 + F23*P31 + F23*P32 + F23*P33 + F23*P34 + F23*P35)*F5 + Q18;

 Pn19 = (F18*P0 + F18*P1 + F18*P2 + F18*P3 + F18*P4 + F18*P5)*F11 + 
    (F19*P6 + F19*P7 + F19*P8 + F19*P9 + F19*P10 + F19*P11)*F11 + 
    (F20*P12 + F20*P13 + F20*P14 + F20*P15 + F20*P16 + F20*P17)*F11 + 
    (F21*P18 + F21*P19 + F21*P20 + F21*P21 + F21*P22 + F21*P23)*F11 + 
    (F22*P24 + F22*P25 + F22*P26 + F22*P27 + F22*P28 + F22*P29)*F11 + 
    (F23*P30 + F23*P31 + F23*P32 + F23*P33 + F23*P34 + F23*P35)*F11 + Q19;

 Pn20 = (F18*P0 + F18*P1 + F18*P2 + F18*P3 + F18*P4 + F18*P5)*F17 + 
    (F19*P6 + F19*P7 + F19*P8 + F19*P9 + F19*P10 + F19*P11)*F17 + 
    (F20*P12 + F20*P13 + F20*P14 + F20*P15 + F20*P16 + F20*P17)*F17 + 
    (F21*P18 + F21*P19 + F21*P20 + F21*P21 + F21*P22 + F21*P23)*F17 + 
    (F22*P24 + F22*P25 + F22*P26 + F22*P27 + F22*P28 + F22*P29)*F17 + 
    (F23*P30 + F23*P31 + F23*P32 + F23*P33 + F23*P34 + F23*P35)*F17 + Q20;

 Pn21 = (F18*P0 + F18*P1 + F18*P2 + F18*P3 + F18*P4 + F18*P5)*F23 + 
    (F19*P6 + F19*P7 + F19*P8 + F19*P9 + F19*P10 + F19*P11)*F23 + 
    (F20*P12 + F20*P13 + F20*P14 + F20*P15 + F20*P16 + F20*P17)*F23 + 
    (F21*P18 + F21*P19 + F21*P20 + F21*P21 + F21*P22 + F21*P23)*F23 + 
    (F22*P24 + F22*P25 + F22*P26 + F22*P27 + F22*P28 + F22*P29)*F23 + 
    (F23*P30 + F23*P31 + F23*P32 + F23*P33 + F23*P34 + F23*P35)*F23 + Q21;

 Pn22 = (F18*P0 + F18*P1 + F18*P2 + F18*P3 + F18*P4 + F18*P5)*F29 + 
    (F19*P6 + F19*P7 + F19*P8 + F19*P9 + F19*P10 + F19*P11)*F29 + 
    (F20*P12 + F20*P13 + F20*P14 + F20*P15 + F20*P16 + F20*P17)*F29 + 
    (F21*P18 + F21*P19 + F21*P20 + F21*P21 + F21*P22 + F21*P23)*F29 + 
    (F22*P24 + F22*P25 + F22*P26 + F22*P27 + F22*P28 + F22*P29)*F29 + 
    (F23*P30 + F23*P31 + F23*P32 + F23*P33 + F23*P34 + F23*P35)*F29 + Q22;

 Pn23 = (F18*P0 + F18*P1 + F18*P2 + F18*P3 + F18*P4 + F18*P5)*F35 + 
    (F19*P6 + F19*P7 + F19*P8 + F19*P9 + F19*P10 + F19*P11)*F35 + 
    (F20*P12 + F20*P13 + F20*P14 + F20*P15 + F20*P16 + F20*P17)*F35 + 
    (F21*P18 + F21*P19 + F21*P20 + F21*P21 + F21*P22 + F21*P23)*F35 + 
    (F22*P24 + F22*P25 + F22*P26 + F22*P27 + F22*P28 + F22*P29)*F35 + 
    (F23*P30 + F23*P31 + F23*P32 + F23*P33 + F23*P34 + F23*P35)*F35 + Q23;

 Pn24 = (F24*P0 + F24*P1 + F24*P2 + F24*P3 + F24*P4 + F24*P5)*F5 + 
    (F25*P6 + F25*P7 + F25*P8 + F25*P9 + F25*P10 + F25*P11)*F5 + 
    (F26*P12 + F26*P13 + F26*P14 + F26*P15 + F26*P16 + F26*P17)*F5 + 
    (F27*P18 + F27*P19 + F27*P20 + F27*P21 + F27*P22 + F27*P23)*F5 + 
    (F28*P24 + F28*P25 + F28*P26 + F28*P27 + F28*P28 + F28*P29)*F5 + 
    (F29*P30 + F29*P31 + F29*P32 + F29*P33 + F29*P34 + F29*P35)*F5 + Q24;

 Pn25 = (F24*P0 + F24*P1 + F24*P2 + F24*P3 + F24*P4 + F24*P5)*F11 + 
    (F25*P6 + F25*P7 + F25*P8 + F25*P9 + F25*P10 + F25*P11)*F11 + 
    (F26*P12 + F26*P13 + F26*P14 + F26*P15 + F26*P16 + F26*P17)*F11 + 
    (F27*P18 + F27*P19 + F27*P20 + F27*P21 + F27*P22 + F27*P23)*F11 + 
    (F28*P24 + F28*P25 + F28*P26 + F28*P27 + F28*P28 + F28*P29)*F11 + 
    (F29*P30 + F29*P31 + F29*P32 + F29*P33 + F29*P34 + F29*P35)*F11 + Q25;

 Pn26 = (F24*P0 + F24*P1 + F24*P2 + F24*P3 + F24*P4 + F24*P5)*F17 + 
    (F25*P6 + F25*P7 + F25*P8 + F25*P9 + F25*P10 + F25*P11)*F17 + 
    (F26*P12 + F26*P13 + F26*P14 + F26*P15 + F26*P16 + F26*P17)*F17 + 
    (F27*P18 + F27*P19 + F27*P20 + F27*P21 + F27*P22 + F27*P23)*F17 + 
    (F28*P24 + F28*P25 + F28*P26 + F28*P27 + F28*P28 + F28*P29)*F17 + 
    (F29*P30 + F29*P31 + F29*P32 + F29*P33 + F29*P34 + F29*P35)*F17 + Q26;

 Pn27 = (F24*P0 + F24*P1 + F24*P2 + F24*P3 + F24*P4 + F24*P5)*F23 + 
    (F25*P6 + F25*P7 + F25*P8 + F25*P9 + F25*P10 + F25*P11)*F23 + 
    (F26*P12 + F26*P13 + F26*P14 + F26*P15 + F26*P16 + F26*P17)*F23 + 
    (F27*P18 + F27*P19 + F27*P20 + F27*P21 + F27*P22 + F27*P23)*F23 + 
    (F28*P24 + F28*P25 + F28*P26 + F28*P27 + F28*P28 + F28*P29)*F23 + 
    (F29*P30 + F29*P31 + F29*P32 + F29*P33 + F29*P34 + F29*P35)*F23 + Q27;

 Pn28 = (F24*P0 + F24*P1 + F24*P2 + F24*P3 + F24*P4 + F24*P5)*F29 + 
    (F25*P6 + F25*P7 + F25*P8 + F25*P9 + F25*P10 + F25*P11)*F29 + 
    (F26*P12 + F26*P13 + F26*P14 + F26*P15 + F26*P16 + F26*P17)*F29 + 
    (F27*P18 + F27*P19 + F27*P20 + F27*P21 + F27*P22 + F27*P23)*F29 + 
    (F28*P24 + F28*P25 + F28*P26 + F28*P27 + F28*P28 + F28*P29)*F29 + 
    (F29*P30 + F29*P31 + F29*P32 + F29*P33 + F29*P34 + F29*P35)*F29 + Q28;

 Pn29 = (F24*P0 + F24*P1 + F24*P2 + F24*P3 + F24*P4 + F24*P5)*F35 + 
    (F25*P6 + F25*P7 + F25*P8 + F25*P9 + F25*P10 + F25*P11)*F35 + 
    (F26*P12 + F26*P13 + F26*P14 + F26*P15 + F26*P16 + F26*P17)*F35 + 
    (F27*P18 + F27*P19 + F27*P20 + F27*P21 + F27*P22 + F27*P23)*F35 + 
    (F28*P24 + F28*P25 + F28*P26 + F28*P27 + F28*P28 + F28*P29)*F35 + 
    (F29*P30 + F29*P31 + F29*P32 + F29*P33 + F29*P34 + F29*P35)*F35 + Q29;

 Pn30 = (F30*P0 + F30*P1 + F30*P2 + F30*P3 + F30*P4 + F30*P5)*F5 + 
    (F31*P6 + F31*P7 + F31*P8 + F31*P9 + F31*P10 + F31*P11)*F5 + 
    (F32*P12 + F32*P13 + F32*P14 + F32*P15 + F32*P16 + F32*P17)*F5 + 
    (F33*P18 + F33*P19 + F33*P20 + F33*P21 + F33*P22 + F33*P23)*F5 + 
    (F34*P24 + F34*P25 + F34*P26 + F34*P27 + F34*P28 + F34*P29)*F5 + 
    (F35*P30 + F35*P31 + F35*P32 + F35*P33 + F35*P34 + F35*P35)*F5 + Q30;

 Pn31 = (F30*P0 + F30*P1 + F30*P2 + F30*P3 + F30*P4 + F30*P5)*F11 + 
    (F31*P6 + F31*P7 + F31*P8 + F31*P9 + F31*P10 + F31*P11)*F11 + 
    (F32*P12 + F32*P13 + F32*P14 + F32*P15 + F32*P16 + F32*P17)*F11 + 
    (F33*P18 + F33*P19 + F33*P20 + F33*P21 + F33*P22 + F33*P23)*F11 + 
    (F34*P24 + F34*P25 + F34*P26 + F34*P27 + F34*P28 + F34*P29)*F11 + 
    (F35*P30 + F35*P31 + F35*P32 + F35*P33 + F35*P34 + F35*P35)*F11 + Q31;

 Pn32 = (F30*P0 + F30*P1 + F30*P2 + F30*P3 + F30*P4 + F30*P5)*F17 + 
    (F31*P6 + F31*P7 + F31*P8 + F31*P9 + F31*P10 + F31*P11)*F17 + 
    (F32*P12 + F32*P13 + F32*P14 + F32*P15 + F32*P16 + F32*P17)*F17 + 
    (F33*P18 + F33*P19 + F33*P20 + F33*P21 + F33*P22 + F33*P23)*F17 + 
    (F34*P24 + F34*P25 + F34*P26 + F34*P27 + F34*P28 + F34*P29)*F17 + 
    (F35*P30 + F35*P31 + F35*P32 + F35*P33 + F35*P34 + F35*P35)*F17 + Q32;

 Pn33 = (F30*P0 + F30*P1 + F30*P2 + F30*P3 + F30*P4 + F30*P5)*F23 + 
    (F31*P6 + F31*P7 + F31*P8 + F31*P9 + F31*P10 + F31*P11)*F23 + 
    (F32*P12 + F32*P13 + F32*P14 + F32*P15 + F32*P16 + F32*P17)*F23 + 
    (F33*P18 + F33*P19 + F33*P20 + F33*P21 + F33*P22 + F33*P23)*F23 + 
    (F34*P24 + F34*P25 + F34*P26 + F34*P27 + F34*P28 + F34*P29)*F23 + 
    (F35*P30 + F35*P31 + F35*P32 + F35*P33 + F35*P34 + F35*P35)*F23 + Q33;

 Pn34 = (F30*P0 + F30*P1 + F30*P2 + F30*P3 + F30*P4 + F30*P5)*F29 + 
    (F31*P6 + F31*P7 + F31*P8 + F31*P9 + F31*P10 + F31*P11)*F29 + 
    (F32*P12 + F32*P13 + F32*P14 + F32*P15 + F32*P16 + F32*P17)*F29 + 
    (F33*P18 + F33*P19 + F33*P20 + F33*P21 + F33*P22 + F33*P23)*F29 + 
    (F34*P24 + F34*P25 + F34*P26 + F34*P27 + F34*P28 + F34*P29)*F29 + 
    (F35*P30 + F35*P31 + F35*P32 + F35*P33 + F35*P34 + F35*P35)*F29 + Q34;

 Pn35 = (F30*P0 + F30*P1 + F30*P2 + F30*P3 + F30*P4 + F30*P5)*F35 + 
    (F31*P6 + F31*P7 + F31*P8 + F31*P9 + F31*P10 + F31*P11)*F35 + 
    (F32*P12 + F32*P13 + F32*P14 + F32*P15 + F32*P16 + F32*P17)*F35 + 
    (F33*P18 + F33*P19 + F33*P20 + F33*P21 + F33*P22 + F33*P23)*F35 + 
    (F34*P24 + F34*P25 + F34*P26 + F34*P27 + F34*P28 + F34*P29)*F35 + 
    (F35*P30 + F35*P31 + F35*P32 + F35*P33 + F35*P34 + F35*P35)*F35 + Q35;
    end
endmodule

`timescale 1ns / 1ps

module Fusion_Unit_tb;

    reg signed [15:0] P1_0,  P1_6,  P1_14, P1_21, P1_28, P1_36;
    reg signed [15:0] P2_0,  P2_6,  P2_14, P2_21, P2_28, P2_36;

    reg signed [15:0] X1_0, X1_1, X1_2, X1_3, X1_4, X1_5;
    reg signed [15:0] X2_0, X2_1, X2_2, X2_3, X2_4, X2_5;

    wire signed [15:0] X0f, X1f, X2f, X3f, X4f, X5f;
    wire signed [31:0] Pf1, Pf2, Pf3, Pf4, Pf5, Pf6;

    Fusion_unit dut (
        .P1_0(P1_0),   .P2_0(P2_0),
        .P1_6(P1_6),   .P2_6(P2_6),
        .P1_14(P1_14), .P2_14(P2_14),
        .P1_21(P1_21), .P2_21(P2_21),
        .P1_28(P1_28), .P2_28(P2_28),
        .P1_36(P1_36), .P2_36(P2_36),

        .X1_0(X1_0), .X2_0(X2_0),
        .X1_1(X1_1), .X2_1(X2_1),
        .X1_2(X1_2), .X2_2(X2_2),
        .X1_3(X1_3), .X2_3(X2_3),
        .X1_4(X1_4), .X2_4(X2_4),
        .X1_5(X1_5), .X2_5(X2_5),

        .X0f(X0f), .X1f(X1f), .X2f(X2f),
        .X3f(X3f), .X4f(X4f), .X5f(X5f),

        .Pf1(Pf1), .Pf2(Pf2), .Pf3(Pf3),
        .Pf4(Pf4), .Pf5(Pf5), .Pf6(Pf6)
    );

    initial begin
        P1_0=0;  P1_6=0;  P1_14=0; P1_21=0; P1_28=0; P1_36=0;
        P2_0=0;  P2_6=0;  P2_14=0; P2_21=0; P2_28=0; P2_36=0;

        X1_0=0; X1_1=0; X1_2=0; X1_3=0; X1_4=0; X1_5=0;
        X2_0=0; X2_1=0; X2_2=0; X2_3=0; X2_4=0; X2_5=0;

        #5;
        P1_0  = 16'd12; P1_6  = 16'd13; P1_14 = 16'd14;
        P1_21 = 16'd15; P1_28 = 16'd16; P1_36 = 16'd17;

        P2_0  = 16'd17; P2_6  = 16'd16; P2_14 = 16'd15;
        P2_21 = 16'd14; P2_28 = 16'd13; P2_36 = 16'd12;

        #5;
        X1_0 = 16'd4; X1_1 = 16'd5; X1_2 = 16'd6;
        X1_3 = 16'd7; X1_4 = 16'd8; X1_5 = 16'd9;

        X2_0 = 16'd9; X2_1 = 16'd8; X2_2 = 16'd7;
        X2_3 = 16'd6; X2_4 = 16'd5; X2_5 = 16'd4;

        #70;
        $finish;
    end

endmodule
